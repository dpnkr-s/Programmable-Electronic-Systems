

  subtype datatype is integer range -65536 to 65535;
  type ioarray is array (0 to 84) of datatype;

  type rom is array (0 to 16) of datatype;
  constant coeff : rom := (-282,
                           -369,
                           -307,
                           -67,
                           326,
                           803,
                           1259,
                           1587,
                           1706,
                           1587,
                           1259,
                           803,
                           326,
                           -67,
                           -307,
                           -369,
                           -282
                           );


  constant inputdata : ioarray := (0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  1,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  0,
                                  -6754,
                                  -15687,
                                  -31716,
                                  -6518,
                                  7301,
                                  -10850,
                                  31710,
                                  -2341,
                                  999,
                                  -30678,
                                  24927,
                                  6725,
                                  -12612,
                                  -7333,
                                  2755,
                                  25075,
                                  24101,
                                  -7305,
                                  10859,
                                  26998,
                                  26665,
                                  152,
                                  -6149,
                                  -17218,
                                  -7584,
                                  16591,
                                  -31878,
                                  32457,
                                  23096,
                                  26618,
                                  27595,
                                  -16927,
                                  -16990,
                                  29897,
                                  24311,
                                  -3735,
                                  -10177,
                                  23941,
                                  -16392,
                                  -11137,
                                  29304,
                                  -5486,
                                  19224,
                                  12300,
                                  -28414,
                                  -24613,
                                  -18685,
                                  11771,
                                  -13118,
                                  -7813,
                                  -25070);

